module DataSyncLib(input clk_100M,input n_rst);



endmodule
